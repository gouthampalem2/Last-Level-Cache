initial 
begin
if($value$plusargs
